module adder32(result, a, b);
   input[31:0] a;
   input[31:0] b;
   output [31:0] result;
   wire [32:0] sum = {1'b0,a} + {1'b0,b};
   assign result = sum[32] ? sum[32:1]: sum[31:0];

endmodule