module cpu( input [31:0] instruction);

endmodule